../ha/ha.sv